module not (
    input wire a,
    output wire q,
) (
    assign q = !a;
);
    
endmodule